`timescale 1ns/1ps
`define T_CLK * 10

module testbench();

wire in_b;
wire in_a;


endmodule